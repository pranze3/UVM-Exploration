package gcd_env_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import gcd_seq_pkg::*;
  import gcd_agent_pkg::*;
  `include "gcd_sb.sv"
  `include "gcd_env.sv"

endpackage : gcd_env_pkg
