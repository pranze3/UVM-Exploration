package gcd_test_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import gcd_env_pkg::*;
  import gcd_seq_pkg::*;
  `include "gcd_base_test.svh"
  `include "gcd_test_lib.sv"
  
endpackage : gcd_test_pkg
