package gcd_seq_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "gcd_seq_item.sv"
  `include "gcd_sequence.svh"
  `include "gcd_seq_lib.sv"
  
endpackage : gcd_seq_pkg
